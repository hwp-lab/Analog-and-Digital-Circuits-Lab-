`timescale 1ns / 1ps
module 7_Segment_Decoder(
    input       [3:0] d,
    output reg  [6:0] cn//cn表示低电平有效，七段字形a, b, … g依次对应y[6], y[5], … y[0]
    );

    always @(*) begin
        case(d)
            4'b0000: cn=7'b00_00001;//0
            4'b0001: cn=7'b100_1111;//1
            4'b0010: cn=7'b001_0010;//2
            4'b0011: cn=7'b000_0110;//3
            4'b0100: cn=7'b100_1100;//4
            4'b0101: cn=7'b010_0100;//5
            4'b0110: cn=7'b010_0000;//6
            4'b0111: cn=7'b000_1111;//7
            4'b1000: cn=7'b000_0000;//8
            4'b1001: cn=7'b000_0100;//9
            4'b1010: cn=7'b000_1000;//a
            4'b1011: cn=7'b110_0000;//b
            4'b1100: cn=7'b011_0001;//c
            4'b1101: cn=7'b100_0010;//d
            4'b1110: cn=7'b011_0000;//e
            4'b1111: cn=7'b011_1000;//f
            default: cn=7'b111_1111;
    endcase
    end
endmodule
