`timescale 1ns / 1ps

module tb_SSD;

    // 输入信号
    reg [3:0] d;
    
    // 输出信号
    wire [6:0] yn;
    
    // 实例化被测试模块
    SSD uut (
        .d(d),
        .yn(yn)
    );
    
    // 测试逻辑
    initial begin
        // 初始化输入
        d = 4'b0000;
        
        // 测试所有BCD输入 (0-9)
        #10 d = 4'b0000; // 0
        #10 d = 4'b0001; // 1
        #10 d = 4'b0010; // 2
        #10 d = 4'b0011; // 3
        #10 d = 4'b0100; // 4
        #10 d = 4'b0101; // 5
        #10 d = 4'b0110; // 6
        #10 d = 4'b0111; // 7
        #10 d = 4'b1000; // 8
        #10 d = 4'b1001; // 9
        
        // 测试非法输入 (10-15)
        #10 d = 4'b1010; // 10
        #10 d = 4'b1011; // 11
        #10 d = 4'b1100; // 12
        #10 d = 4'b1101; // 13
        #10 d = 4'b1110; // 14
        #10 d = 4'b1111; // 15
        
        #10 $finish;
    end
endmodule